package UART_PACKAGE; 
    parameter DATA_WIDTH = 8;
endpackage : UART_PACKAGE 